`include "components/alu.v"
`include "components/adder.v"
`include "components/datamemory.v"
`include "components/instructiondecode.v"
`include "components/muxes.v"
`include "components/pc.v"
`include "components/regfile.v"
`include "components/shifter.v"
`include "components/signextend.v"


module cpu();

endmodule