`include "components/alu.v"

module cpu();

endmodule